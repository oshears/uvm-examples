`timescale 1ns/1ns
package GamePackage;

    localparam int NUM_ROWS = 6;
    localparam int NUM_COLS = 7;

endpackage : GamePackage
