`timescale 1ns/1ns
package GamePackage;

    const int NUM_ROWS = 6;
    const int NUM_COLS = 7;

endpackage : GamePackage
