`timescale 1ns/1ns
class Board;

    // OYS: Use unpacked array because the data is all independent
    // Columns x Rows
    int board[7][6];

    string boardName;

    // static const NUM_ROWS

    // static const int NUM_ROWS = 6;
    // static const int NUM_COLS = 7;

    function new (string boardName = "Default Board");
        this.boardName = boardName;
        // no need to initialize board since its statically allocated
    endfunction

    function void PlaceInColumn(int column, int value);
        board[column][0] = value;
    endfunction

    function void PlaceAtPosition(int col, int row, int value);
        board[col][row] = value;
    endfunction

    function int NextEmptySpace(int column); 
    // this func returns the value of row

        foreach (board[column][row]) begin // row is the iterator
            if (row == 0) begin
                return row;
                // alternatively you can set the result to the function name
                // e.g., NextEmptySpace = row
                // you can also declare input/output directions in the function name
                // that would allow you to return multiple values
            end
        end

    endfunction

    function void ResetBoard();
        board = '{default: 0};
    endfunction

    function void Display();

        for(int row = 5; row > -1; row--) begin
            for(int col = 0; col < 7; col++) begin
                $write("%d",board[col][row]);
            end
            $display("");
        end
    endfunction


endclass